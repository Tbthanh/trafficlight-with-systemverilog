module trafficlight (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	input car,

	output light
);

	
endmodule : trafficlight